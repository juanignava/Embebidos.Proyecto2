// sistema_tb.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module sistema_tb (
	);

	wire        sistema_inst_clk_bfm_clk_clk;       // sistema_inst_clk_bfm:clk -> [sistema_inst:clk_clk, sistema_inst_reset_bfm:clk]
	wire  [7:0] sistema_inst_regs_export;           // sistema_inst:regs_export -> sistema_inst_regs_bfm:sig_export
	wire        sistema_inst_reset_bfm_reset_reset; // sistema_inst_reset_bfm:reset -> sistema_inst:reset_reset_n

	sistema sistema_inst (
		.clk_clk       (sistema_inst_clk_bfm_clk_clk),       //   clk.clk
		.regs_export   (sistema_inst_regs_export),           //  regs.export
		.reset_reset_n (sistema_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sistema_inst_clk_bfm (
		.clk (sistema_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm sistema_inst_regs_bfm (
		.sig_export (sistema_inst_regs_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sistema_inst_reset_bfm (
		.reset (sistema_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sistema_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
