// alarm_clk_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module alarm_clk_tb (
	);

	wire        alarm_clk_inst_clk_bfm_clk_clk;                 // alarm_clk_inst_clk_bfm:clk -> [alarm_clk_inst:clk_clk, alarm_clk_inst_reset_bfm:clk]
	wire        alarm_clk_inst_alarm_export;                    // alarm_clk_inst:alarm_export -> alarm_clk_inst_alarm_bfm:sig_export
	wire  [0:0] alarm_clk_inst_btn_down_bfm_conduit_export;     // alarm_clk_inst_btn_down_bfm:sig_export -> alarm_clk_inst:btn_down_export
	wire  [0:0] alarm_clk_inst_btn_set_bfm_conduit_export;      // alarm_clk_inst_btn_set_bfm:sig_export -> alarm_clk_inst:btn_set_export
	wire  [0:0] alarm_clk_inst_btn_up_bfm_conduit_export;       // alarm_clk_inst_btn_up_bfm:sig_export -> alarm_clk_inst:btn_up_export
	wire  [3:0] alarm_clk_inst_display_h0_export;               // alarm_clk_inst:display_h0_export -> alarm_clk_inst_display_h0_bfm:sig_export
	wire  [3:0] alarm_clk_inst_display_h1_export;               // alarm_clk_inst:display_h1_export -> alarm_clk_inst_display_h1_bfm:sig_export
	wire  [3:0] alarm_clk_inst_display_m0_export;               // alarm_clk_inst:display_m0_export -> alarm_clk_inst_display_m0_bfm:sig_export
	wire  [3:0] alarm_clk_inst_display_m1_export;               // alarm_clk_inst:display_m1_export -> alarm_clk_inst_display_m1_bfm:sig_export
	wire  [3:0] alarm_clk_inst_display_s0_export;               // alarm_clk_inst:display_s0_export -> alarm_clk_inst_display_s0_bfm:sig_export
	wire  [3:0] alarm_clk_inst_display_s1_export;               // alarm_clk_inst:display_s1_export -> alarm_clk_inst_display_s1_bfm:sig_export
	wire  [0:0] alarm_clk_inst_swc_activate_bfm_conduit_export; // alarm_clk_inst_swc_activate_bfm:sig_export -> alarm_clk_inst:swc_activate_export
	wire  [0:0] alarm_clk_inst_swc_sel_bfm_conduit_export;      // alarm_clk_inst_swc_sel_bfm:sig_export -> alarm_clk_inst:swc_sel_export
	wire        alarm_clk_inst_reset_bfm_reset_reset;           // alarm_clk_inst_reset_bfm:reset -> alarm_clk_inst:reset_reset_n

	alarm_clk alarm_clk_inst (
		.alarm_export        (alarm_clk_inst_alarm_export),                    //        alarm.export
		.btn_down_export     (alarm_clk_inst_btn_down_bfm_conduit_export),     //     btn_down.export
		.btn_set_export      (alarm_clk_inst_btn_set_bfm_conduit_export),      //      btn_set.export
		.btn_up_export       (alarm_clk_inst_btn_up_bfm_conduit_export),       //       btn_up.export
		.clk_clk             (alarm_clk_inst_clk_bfm_clk_clk),                 //          clk.clk
		.display_h0_export   (alarm_clk_inst_display_h0_export),               //   display_h0.export
		.display_h1_export   (alarm_clk_inst_display_h1_export),               //   display_h1.export
		.display_m0_export   (alarm_clk_inst_display_m0_export),               //   display_m0.export
		.display_m1_export   (alarm_clk_inst_display_m1_export),               //   display_m1.export
		.display_s0_export   (alarm_clk_inst_display_s0_export),               //   display_s0.export
		.display_s1_export   (alarm_clk_inst_display_s1_export),               //   display_s1.export
		.reset_reset_n       (alarm_clk_inst_reset_bfm_reset_reset),           //        reset.reset_n
		.swc_activate_export (alarm_clk_inst_swc_activate_bfm_conduit_export), // swc_activate.export
		.swc_sel_export      (alarm_clk_inst_swc_sel_bfm_conduit_export)       //      swc_sel.export
	);

	altera_conduit_bfm alarm_clk_inst_alarm_bfm (
		.sig_export (alarm_clk_inst_alarm_export)  // conduit.export
	);

	altera_conduit_bfm_0002 alarm_clk_inst_btn_down_bfm (
		.sig_export (alarm_clk_inst_btn_down_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 alarm_clk_inst_btn_set_bfm (
		.sig_export (alarm_clk_inst_btn_set_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 alarm_clk_inst_btn_up_bfm (
		.sig_export (alarm_clk_inst_btn_up_bfm_conduit_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) alarm_clk_inst_clk_bfm (
		.clk (alarm_clk_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0003 alarm_clk_inst_display_h0_bfm (
		.sig_export (alarm_clk_inst_display_h0_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarm_clk_inst_display_h1_bfm (
		.sig_export (alarm_clk_inst_display_h1_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarm_clk_inst_display_m0_bfm (
		.sig_export (alarm_clk_inst_display_m0_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarm_clk_inst_display_m1_bfm (
		.sig_export (alarm_clk_inst_display_m1_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarm_clk_inst_display_s0_bfm (
		.sig_export (alarm_clk_inst_display_s0_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarm_clk_inst_display_s1_bfm (
		.sig_export (alarm_clk_inst_display_s1_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) alarm_clk_inst_reset_bfm (
		.reset (alarm_clk_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (alarm_clk_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 alarm_clk_inst_swc_activate_bfm (
		.sig_export (alarm_clk_inst_swc_activate_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 alarm_clk_inst_swc_sel_bfm (
		.sig_export (alarm_clk_inst_swc_sel_bfm_conduit_export)  // conduit.export
	);

endmodule
